// Copyright 2021 OpenHW Group
// Copyright 2021 Datum Technology Corporation
// Copyright 2021 Silicon Labs
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_MEM_CONSTANTS_SV__
`define __UVML_MEM_CONSTANTS_SV__




`endif // __UVML_MEM_CONSTANTS_SV__
