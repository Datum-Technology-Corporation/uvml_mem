// Copyright 2021 OpenHW Group
// Copyright 2021 Datum Technology Corporation
// Copyright 2021 Silicon Labs
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_MEM_MACROS_SV__
`define __UVML_MEM_MACROS_SV__


`define UVML_MEM_DEFAULT_XLEN   32
`define UVML_MEM_DEFAULT_NBYTES  4


`endif // __UVML_MEM_MACROS_SV__
